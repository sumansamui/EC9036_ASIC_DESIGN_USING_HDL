LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY counter2_tb IS
END counter2_tb;
 
ARCHITECTURE behavior OF counter_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT counter
    PORT(
         clk : IN  std_logic;
         reset : IN  std_logic;
         count : OUT  std_logic_vector(3 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic;
   signal reset : std_logic;

 	--Outputs
   signal count : std_logic_vector(3 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: counter2 PORT MAP (clk => clk, reset => reset, count => count);

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process of reset signal
   stim_proc: process
   begin		
		
		reset<='1';
      -- hold reset state for 100 ns.
      wait for 100 ns;	

		
		reset<='0';

      wait;
   end process;

END;

`timescale 1ns / 1ps

module counter(
    input clk,
    input rst,
    output reg [3:0] count
    );
always @(posedge clk or posedge rst)
begin  
if(rst)
	count<=4'b0000;
else
   count<=count + 1; 
end
endmodule
